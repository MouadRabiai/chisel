module DeviceUnderTestPrintf(
  input        clock,
  input        reset,
  input  [1:0] io_a,
  input  [1:0] io_b,
  output [1:0] io_out
);
  assign io_out = io_a & io_b; // @[DeviceUnderTestPrintf.scala 21:16]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset) begin
          $fwrite(32'h80000002,"dut: %d %d %d\n",io_a,io_b,io_out); // @[DeviceUnderTestPrintf.scala 22:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
